package pkg;

	import uvm_pkg::*;

	`include "uvm_macros.svh"

	`include "ahb_agt_config.sv"
	`include "apb_agt_config.sv"
	`include "env_config.sv"

	
	`include "ahb_xtn.sv"
	`include "apb_xtn.sv"

	`include "ahb_driver.sv"
	`include "ahb_monitor.sv"
	`include "ahb_sequencer.sv"
	`include "ahb_agent.sv"
	`include "ahb_agt_top.sv"
	`include "ahb_seqs.sv"


	`include "apb_driver.sv"
	`include "apb_monitor.sv"
	`include "apb_sequencer.sv"
	`include "apb_agent.sv"
	`include "apb_agt_top.sv"
	`include "apb_seqs.sv"

	
	
	`include "v_sequencer.sv"
	//`include "v_seqs.sv"
	`include "sb.sv"
	`include "env.sv"
	`include "test.sv"

	
endpackage
